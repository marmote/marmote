library verilog;
use verilog.vl_types.all;
entity F2DSS_COMMSMATRIX is
    port(
        HCLK            : in     vl_logic;
        HRESETn         : in     vl_logic;
        F2_TESTREMAPENABLE: in     vl_logic;
        F2_TESTESRAM1REMAP: in     vl_logic;
        F2_ESRAMSIZE    : in     vl_logic_vector(1 downto 0);
        F2_ENVMPOWEREDDOWN: in     vl_logic;
        COM_ESRAMFWREMAP: in     vl_logic;
        COM_ENVMREMAPSIZE: in     vl_logic_vector(4 downto 0);
        COM_ENVMREMAPBASE: in     vl_logic_vector(19 downto 0);
        COM_ENVMFABREMAPBASE: in     vl_logic_vector(19 downto 0);
        COM_PROTREGIONSIZE: in     vl_logic_vector(4 downto 0);
        COM_PROTREGIONBASE: in     vl_logic_vector(31 downto 0);
        COM_MASTERENABLE: in     vl_logic_vector(2 downto 0);
        COM_CLEARSTATUS : in     vl_logic_vector(4 downto 0);
        COM_WEIGHTEDMODE: in     vl_logic;
        COM_ERRORSTATUS : out    vl_logic_vector(4 downto 0);
        COM_ERRORINTERRUPT: out    vl_logic;
        M3_HADDRI       : in     vl_logic_vector(31 downto 0);
        M3_HTRANSI1     : in     vl_logic;
        M3_HSIZEI       : in     vl_logic_vector(2 downto 0);
        M3_HADDRD       : in     vl_logic_vector(31 downto 0);
        M3_HTRANSD1     : in     vl_logic;
        M3_HWRITED      : in     vl_logic;
        M3_HSIZED       : in     vl_logic_vector(2 downto 0);
        M3_HWDATAD      : in     vl_logic_vector(31 downto 0);
        M3_HRDATAI      : out    vl_logic_vector(31 downto 0);
        M3_HREADYI      : out    vl_logic;
        M3_HRESPI       : out    vl_logic;
        M3_HRDATAD      : out    vl_logic_vector(31 downto 0);
        M3_HREADYD      : out    vl_logic;
        M3_HRESPD       : out    vl_logic;
        M3_HADDRS       : in     vl_logic_vector(31 downto 0);
        M3_HTRANSS1     : in     vl_logic;
        M3_HWRITES      : in     vl_logic;
        M3_HSIZES       : in     vl_logic_vector(2 downto 0);
        M3_HWDATAS      : in     vl_logic_vector(31 downto 0);
        M3_HMASTLOCKS   : in     vl_logic;
        M3_HRDATAS      : out    vl_logic_vector(31 downto 0);
        M3_HREADYS      : out    vl_logic;
        M3_HRESPS       : out    vl_logic;
        DS_FM_HADDR     : in     vl_logic_vector(31 downto 0);
        DS_FM_HMASTLOCK : in     vl_logic;
        DS_FM_HSIZE     : in     vl_logic_vector(2 downto 0);
        DS_FM_HTRANS1   : in     vl_logic;
        DS_FM_HWRITE    : in     vl_logic;
        DS_FM_HWDATA    : in     vl_logic_vector(31 downto 0);
        DS_FM_HRDATA    : out    vl_logic_vector(31 downto 0);
        DS_FM_HREADY    : out    vl_logic;
        DS_FM_HRESP     : out    vl_logic;
        MAC_HWRITE      : in     vl_logic;
        MAC_HADDR       : in     vl_logic_vector(31 downto 0);
        MAC_HTRANS1     : in     vl_logic;
        MAC_HSIZE       : in     vl_logic_vector(2 downto 0);
        MAC_HWDATA      : in     vl_logic_vector(31 downto 0);
        MAC_HRDATA      : out    vl_logic_vector(31 downto 0);
        MAC_HREADY      : out    vl_logic;
        MAC_HRESP       : out    vl_logic;
        PDMA_HADDR      : in     vl_logic_vector(31 downto 0);
        PDMA_HSIZE      : in     vl_logic_vector(2 downto 0);
        PDMA_HTRANS1    : in     vl_logic;
        PDMA_HWDATA     : in     vl_logic_vector(31 downto 0);
        PDMA_HWRITE     : in     vl_logic;
        PDMA_HRDATA     : out    vl_logic_vector(31 downto 0);
        PDMA_HREADY     : out    vl_logic;
        PDMA_HRESP      : out    vl_logic;
        ESRAM0_HRDATA   : in     vl_logic_vector(31 downto 0);
        ESRAM0_HREADYOUT: in     vl_logic;
        ESRAM0_HRESP    : in     vl_logic;
        ESRAM0_HADDR    : out    vl_logic_vector(31 downto 0);
        ESRAM0_HSIZE    : out    vl_logic_vector(2 downto 0);
        ESRAM0_HTRANS1  : out    vl_logic;
        ESRAM0_HWDATA   : out    vl_logic_vector(31 downto 0);
        ESRAM0_HWRITE   : out    vl_logic;
        ESRAM0_HSEL     : out    vl_logic;
        ESRAM0_HREADY   : out    vl_logic;
        ESRAM1_HRDATA   : in     vl_logic_vector(31 downto 0);
        ESRAM1_HREADYOUT: in     vl_logic;
        ESRAM1_HRESP    : in     vl_logic;
        ESRAM1_HADDR    : out    vl_logic_vector(31 downto 0);
        ESRAM1_HSIZE    : out    vl_logic_vector(2 downto 0);
        ESRAM1_HTRANS1  : out    vl_logic;
        ESRAM1_HWDATA   : out    vl_logic_vector(31 downto 0);
        ESRAM1_HWRITE   : out    vl_logic;
        ESRAM1_HSEL     : out    vl_logic;
        ESRAM1_HREADY   : out    vl_logic;
        ENVM_HRDATA     : in     vl_logic_vector(31 downto 0);
        ENVM_HREADYOUT  : in     vl_logic;
        ENVM_HRESP      : in     vl_logic;
        ENVM_HADDR      : out    vl_logic_vector(31 downto 0);
        ENVM_HSIZE      : out    vl_logic_vector(2 downto 0);
        ENVM_HTRANS1    : out    vl_logic;
        ENVM_HWDATA     : out    vl_logic_vector(31 downto 0);
        ENVM_HWRITE     : out    vl_logic;
        ENVM_HSEL       : out    vl_logic;
        ENVM_HREADY     : out    vl_logic;
        EM_HRDATA       : in     vl_logic_vector(31 downto 0);
        EM_HREADYOUT    : in     vl_logic;
        EM_HRESP        : in     vl_logic;
        EM_HADDR        : out    vl_logic_vector(31 downto 0);
        EM_HSIZE        : out    vl_logic_vector(2 downto 0);
        EM_HTRANS1      : out    vl_logic;
        EM_HWDATA       : out    vl_logic_vector(31 downto 0);
        EM_HWRITE       : out    vl_logic;
        EM_HSEL         : out    vl_logic;
        EM_HREADY       : out    vl_logic;
        ACE_HRDATA      : in     vl_logic_vector(31 downto 0);
        ACE_HREADYOUT   : in     vl_logic;
        ACE_HRESP       : in     vl_logic;
        ACE_HADDR       : out    vl_logic_vector(31 downto 0);
        ACE_HSIZE       : out    vl_logic_vector(2 downto 0);
        ACE_HTRANS1     : out    vl_logic;
        ACE_HREADY      : out    vl_logic;
        ACE_HWDATA      : out    vl_logic_vector(31 downto 0);
        ACE_HWRITE      : out    vl_logic;
        ACE_HSEL        : out    vl_logic;
        DS_HM_HRDATA    : in     vl_logic_vector(31 downto 0);
        DS_HM_HREADYOUT : in     vl_logic;
        DS_HM_HRESP     : in     vl_logic;
        DS_HM_HADDR     : out    vl_logic_vector(31 downto 0);
        DS_HM_HSIZE     : out    vl_logic_vector(2 downto 0);
        DS_HM_HTRANS1   : out    vl_logic;
        DS_HM_HSEL      : out    vl_logic;
        DS_HM_HWRITE    : out    vl_logic;
        DS_HM_HWDATA    : out    vl_logic_vector(31 downto 0);
        DS_HM_HREADY    : out    vl_logic;
        DS_HM_HMASTLOCK : out    vl_logic;
        PER0_HRDATA     : in     vl_logic_vector(31 downto 0);
        PER0_HREADYOUT  : in     vl_logic;
        PER0_HRESP      : in     vl_logic;
        PER0_HADDR      : out    vl_logic_vector(31 downto 0);
        PER0_HSIZE      : out    vl_logic_vector(2 downto 0);
        PER0_HTRANS1    : out    vl_logic;
        PER0_HREADY     : out    vl_logic;
        PER0_HWDATA     : out    vl_logic_vector(31 downto 0);
        PER0_HWRITE     : out    vl_logic;
        PER0_HSEL       : out    vl_logic;
        PER1_HRDATA     : in     vl_logic_vector(31 downto 0);
        PER1_HREADYOUT  : in     vl_logic;
        PER1_HRESP      : in     vl_logic;
        PER1_HADDR      : out    vl_logic_vector(31 downto 0);
        PER1_HSIZE      : out    vl_logic_vector(2 downto 0);
        PER1_HTRANS1    : out    vl_logic;
        PER1_HREADY     : out    vl_logic;
        PER1_HWDATA     : out    vl_logic_vector(31 downto 0);
        PER1_HWRITE     : out    vl_logic;
        PER1_HSEL       : out    vl_logic
    );
end F2DSS_COMMSMATRIX;
