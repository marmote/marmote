library verilog;
use verilog.vl_types.all;
entity F2DSS_FABRICIF is
    port(
        F2_LARGE_CT_XS  : in     vl_logic;
        FPGAGOOD        : in     vl_logic;
        FAB_AHBIF       : in     vl_logic;
        FAB_APB32       : in     vl_logic;
        GLBDIVISOR      : in     vl_logic_vector(1 downto 0);
        FAB_AHB_BYPASS  : in     vl_logic;
        F2_INTCLK       : in     vl_logic;
        APB16_XHOLD     : out    vl_logic_vector(15 downto 0);
        DS_HCLK         : in     vl_logic;
        DS_HRESETN      : in     vl_logic;
        DS_HM_HADDR     : in     vl_logic_vector(19 downto 0);
        DS_HM_HMASTLOCK : in     vl_logic;
        DS_HM_HSIZE     : in     vl_logic_vector(1 downto 0);
        DS_HM_HTRANS1   : in     vl_logic;
        DS_HM_HSEL      : in     vl_logic;
        DS_HM_HWRITE    : in     vl_logic;
        DS_HM_HWDATA    : in     vl_logic_vector(31 downto 0);
        DS_HM_HREADY    : in     vl_logic;
        DS_HM_HREADYOUT : out    vl_logic;
        DS_HM_HRESP     : out    vl_logic;
        DS_HM_HRDATA    : out    vl_logic_vector(31 downto 0);
        F_HM_ADDR       : out    vl_logic_vector(19 downto 0);
        F_HM_WDATA      : out    vl_logic_vector(31 downto 0);
        F_HM_RDATA      : in     vl_logic_vector(31 downto 0);
        F_HM_HMASTLOCK  : out    vl_logic;
        F_HM_HSIZE      : out    vl_logic_vector(1 downto 0);
        F_HM_HTRANS1    : out    vl_logic;
        F_HM_HWRITE     : out    vl_logic;
        F_HM_HREADY     : in     vl_logic;
        F_HM_HRESP      : in     vl_logic;
        F_HM_PSEL       : out    vl_logic;
        F_HM_PENABLE    : out    vl_logic;
        F_HM_PWRITE     : out    vl_logic;
        F_HM_PREADY     : in     vl_logic;
        F_HM_PSLVERR    : in     vl_logic;
        DS_FM_HADDR     : out    vl_logic_vector(31 downto 0);
        DS_FM_HMASTLOCK : out    vl_logic;
        DS_FM_HSIZE     : out    vl_logic_vector(1 downto 0);
        DS_FM_HTRANS1   : out    vl_logic;
        DS_FM_HWRITE    : out    vl_logic;
        DS_FM_HWDATA    : out    vl_logic_vector(31 downto 0);
        DS_FM_HRDATA    : in     vl_logic_vector(31 downto 0);
        DS_FM_HREADY    : in     vl_logic;
        DS_FM_HRESP     : in     vl_logic;
        F_FM_ADDR       : in     vl_logic_vector(31 downto 0);
        F_FM_WDATA      : in     vl_logic_vector(31 downto 0);
        F_FM_RDATA      : out    vl_logic_vector(31 downto 0);
        F_FM_HMASTLOCK  : in     vl_logic;
        F_FM_HSIZE      : in     vl_logic_vector(1 downto 0);
        F_FM_HTRANS1    : in     vl_logic;
        F_FM_HSEL       : in     vl_logic;
        F_FM_HWRITE     : in     vl_logic;
        F_FM_HREADY     : in     vl_logic;
        F_FM_HREADYOUT  : out    vl_logic;
        F_FM_HRESP      : out    vl_logic;
        F_FM_PSEL       : in     vl_logic;
        F_FM_PENABLE    : in     vl_logic;
        F_FM_PWRITE     : in     vl_logic;
        F_FM_PREADY     : out    vl_logic;
        F_FM_PSLVERR    : out    vl_logic;
        CALIBSTART      : in     vl_logic;
        CALIBFAIL       : out    vl_logic;
        F2HCALIB        : in     vl_logic;
        H2FCALIB        : out    vl_logic
    );
end F2DSS_FABRICIF;
