library verilog;
use verilog.vl_types.all;
entity CMSlaveStage is
    port(
        HCLK            : in     vl_logic;
        HRESETn         : in     vl_logic;
        HREADYOUT       : in     vl_logic;
        HRESP           : in     vl_logic;
        HSEL            : out    vl_logic;
        HADDR           : out    vl_logic_vector(31 downto 0);
        HSIZE           : out    vl_logic_vector(2 downto 0);
        HTRANS1         : out    vl_logic;
        HWRITE          : out    vl_logic;
        HWDATA          : out    vl_logic_vector(31 downto 0);
        HREADY_S        : out    vl_logic;
        HMASTLOCK       : out    vl_logic;
        COM_WEIGHTEDMODE: in     vl_logic;
        mAddrSel        : in     vl_logic_vector(4 downto 0);
        mDataSel        : in     vl_logic_vector(4 downto 0);
        mPrevDataSlaveReady: in     vl_logic_vector(4 downto 0);
        mAddrReady      : out    vl_logic_vector(4 downto 0);
        mDataReady      : out    vl_logic_vector(4 downto 0);
        mHResp          : out    vl_logic_vector(4 downto 0);
        m0GatedHADDR    : in     vl_logic_vector(31 downto 0);
        m0GatedHMASTLOCK: in     vl_logic;
        m0GatedHSIZE    : in     vl_logic_vector(2 downto 0);
        m0GatedHTRANS1  : in     vl_logic;
        m0GatedHWRITE   : in     vl_logic;
        m1GatedHADDR    : in     vl_logic_vector(31 downto 0);
        m1GatedHMASTLOCK: in     vl_logic;
        m1GatedHSIZE    : in     vl_logic_vector(2 downto 0);
        m1GatedHTRANS1  : in     vl_logic;
        m1GatedHWRITE   : in     vl_logic;
        m2GatedHADDR    : in     vl_logic_vector(31 downto 0);
        m2GatedHMASTLOCK: in     vl_logic;
        m2GatedHSIZE    : in     vl_logic_vector(2 downto 0);
        m2GatedHTRANS1  : in     vl_logic;
        m2GatedHWRITE   : in     vl_logic;
        m3GatedHADDR    : in     vl_logic_vector(31 downto 0);
        m3GatedHMASTLOCK: in     vl_logic;
        m3GatedHSIZE    : in     vl_logic_vector(2 downto 0);
        m3GatedHTRANS1  : in     vl_logic;
        m3GatedHWRITE   : in     vl_logic;
        m4GatedHADDR    : in     vl_logic_vector(31 downto 0);
        m4GatedHMASTLOCK: in     vl_logic;
        m4GatedHSIZE    : in     vl_logic_vector(2 downto 0);
        m4GatedHTRANS1  : in     vl_logic;
        m4GatedHWRITE   : in     vl_logic;
        HWDATA_M0       : in     vl_logic_vector(31 downto 0);
        HWDATA_M1       : in     vl_logic_vector(31 downto 0);
        HWDATA_M2       : in     vl_logic_vector(31 downto 0);
        HWDATA_M3       : in     vl_logic_vector(31 downto 0);
        HWDATA_M4       : in     vl_logic_vector(31 downto 0)
    );
end CMSlaveStage;
