library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_PPE_RDMUX is
    port(
        RAM_RD_B_apbrd_pre: in     vl_logic;
        RAM_DO_B        : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_CTRL  : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_STATUS: in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA  : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA_PEEK: in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA0 : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA1 : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA2 : in     vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA3 : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_CTRL  : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_STATUS: in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA  : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA_PEEK: in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA0 : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA1 : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA2 : in     vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA3 : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_CTRL  : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_STATUS: in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA  : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA_PEEK: in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA0 : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA1 : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA2 : in     vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA3 : in     vl_logic_vector(31 downto 0);
        PPE_CTRL        : in     vl_logic_vector(31 downto 0);
        PPE_PC_ETC      : in     vl_logic_vector(31 downto 0);
        PPE_SCRATCH     : in     vl_logic_vector(31 downto 0);
        PPE_SF          : in     vl_logic_vector(31 downto 0);
        ALU_CTRL        : in     vl_logic_vector(31 downto 0);
        ALU_STATUS      : in     vl_logic_vector(31 downto 0);
        ALU_A           : in     vl_logic_vector(31 downto 0);
        ALU_B           : in     vl_logic_vector(31 downto 0);
        ALU_C           : in     vl_logic_vector(31 downto 0);
        ALU_D           : in     vl_logic_vector(15 downto 0);
        ALU_E           : in     vl_logic_vector(15 downto 0);
        PPE_FPTR        : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS0      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS1      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS2      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS3      : in     vl_logic_vector(31 downto 0);
        PPE_SFFLAGS     : in     vl_logic_vector(31 downto 0);
        PADDR           : in     vl_logic_vector(12 downto 0);
        PRDATA_PPE      : out    vl_logic_vector(31 downto 0)
    );
end F2DSS_ACE_PPE_RDMUX;
