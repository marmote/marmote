library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_MISC is
    port(
        PCLK            : in     vl_logic;
        PRESETN         : in     vl_logic;
        PADDR           : in     vl_logic_vector(12 downto 0);
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PRDATA_SSE      : in     vl_logic_vector(15 downto 0);
        PRDATA_PPE      : in     vl_logic_vector(31 downto 0);
        PREADY_SSE      : in     vl_logic;
        PREADY_PPE      : in     vl_logic;
        PSEL_SSE        : out    vl_logic;
        PSEL_PPE        : out    vl_logic;
        PRDATA          : out    vl_logic_vector(31 downto 0);
        PREADY          : out    vl_logic;
        PSLVERR         : out    vl_logic;
        PPE_PDMA_DATAOUT_reg_move_target: in     vl_logic;
        PPE_PDMA_DATAOUT_chan_en: in     vl_logic;
        PPE_PDMA_DATAOUT_raw_en: in     vl_logic;
        PPE_PDMA_DATAOUT_tag_en: in     vl_logic;
        PPE_PDMA_CTRL_reg_move_target: in     vl_logic;
        xfer_din_mux    : in     vl_logic_vector(31 downto 0);
        CURRENT_ADC_CHAN: in     vl_logic_vector(5 downto 0);
        ACE_INREADY     : in     vl_logic;
        ACE_OUTREADY    : out    vl_logic;
        ADC0_CALIBRATE  : in     vl_logic;
        ADC1_CALIBRATE  : in     vl_logic;
        ADC2_CALIBRATE  : in     vl_logic;
        ADC0_SAMPLE     : in     vl_logic;
        ADC1_SAMPLE     : in     vl_logic;
        ADC2_SAMPLE     : in     vl_logic;
        ADC0_BUSY       : in     vl_logic;
        ADC1_BUSY       : in     vl_logic;
        ADC2_BUSY       : in     vl_logic;
        ADC0_DATAVALID  : in     vl_logic;
        ADC1_DATAVALID  : in     vl_logic;
        ADC2_DATAVALID  : in     vl_logic;
        ADC0_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC1_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC2_RESULT     : in     vl_logic_vector(11 downto 0);
        COMPARATOR      : in     vl_logic_vector(11 downto 0);
        ADC0_CALIBRATE_rise: in     vl_logic;
        ADC1_CALIBRATE_rise: in     vl_logic;
        ADC2_CALIBRATE_rise: in     vl_logic;
        ADC0_CALIBRATE_fall: in     vl_logic;
        ADC1_CALIBRATE_fall: in     vl_logic;
        ADC2_CALIBRATE_fall: in     vl_logic;
        ADC0_DATAVALID_rise: in     vl_logic;
        ADC1_DATAVALID_rise: in     vl_logic;
        ADC2_DATAVALID_rise: in     vl_logic;
        PC0_FLAGS       : in     vl_logic_vector(3 downto 0);
        PC1_FLAGS       : in     vl_logic_vector(3 downto 0);
        PC2_FLAGS       : in     vl_logic_vector(3 downto 0);
        PPE_FLAGS0      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS1      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS2      : in     vl_logic_vector(31 downto 0);
        PPE_FLAGS3      : in     vl_logic_vector(31 downto 0);
        PPE_SFFLAGS     : in     vl_logic_vector(31 downto 0);
        PPE_BUSY        : in     vl_logic;
        ADC0_FIFO_FULL  : in     vl_logic;
        ADC0_FIFO_AFULL : in     vl_logic;
        ADC1_FIFO_FULL  : in     vl_logic;
        ADC1_FIFO_AFULL : in     vl_logic;
        ADC2_FIFO_FULL  : in     vl_logic;
        ADC2_FIFO_AFULL : in     vl_logic;
        ADC0_FIFO_EMPTY : in     vl_logic;
        ADC1_FIFO_EMPTY : in     vl_logic;
        ADC2_FIFO_EMPTY : in     vl_logic;
        FPGA_FLAGS      : out    vl_logic_vector(31 downto 0);
        INTERRUPT       : out    vl_logic_vector(85 downto 0)
    );
end F2DSS_ACE_MISC;
