library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_PPE_ALU is
    port(
        PCLK            : in     vl_logic;
        PRESETN         : in     vl_logic;
        PADDR           : in     vl_logic_vector(12 downto 0);
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PPE_BUSY        : in     vl_logic;
        CURRENT_ADC_CHAN: in     vl_logic_vector(5 downto 0);
        RAM_DO_A        : in     vl_logic_vector(31 downto 0);
        PC_inc          : in     vl_logic;
        PC_init_addr_ld : in     vl_logic;
        PC_init_addr    : in     vl_logic_vector(9 downto 0);
        PC_ETC_busy     : in     vl_logic;
        SF_busy         : in     vl_logic;
        SCRATCH_busy    : in     vl_logic;
        ALU_CTRL_busy   : in     vl_logic;
        A_busy          : in     vl_logic;
        B_busy          : in     vl_logic;
        C_busy          : in     vl_logic;
        D_busy          : in     vl_logic;
        E_busy          : in     vl_logic;
        Ci_busy         : in     vl_logic;
        NegA_busy       : in     vl_logic;
        C2a_busy        : in     vl_logic;
        s2B_busy        : in     vl_logic;
        C2d_busy        : in     vl_logic;
        st_filt_cnt_clr : in     vl_logic;
        st_filt_cnt_inc : in     vl_logic;
        st_filt_st_one  : in     vl_logic;
        st_filt_st_zero : in     vl_logic;
        PPE_thresh_op_load: in     vl_logic;
        xfer_load_special_active: in     vl_logic;
        xfer_move_active: in     vl_logic;
        PPE_CTRL_reg_move_target: in     vl_logic;
        PC_ETC_reg_move_target: in     vl_logic;
        SCRATCH_reg_move_target: in     vl_logic;
        SF_reg_move_target: in     vl_logic;
        ALU_CTRL_reg_move_target: in     vl_logic;
        A_reg_move_target: in     vl_logic;
        B_reg_move_target: in     vl_logic;
        C_reg_move_target: in     vl_logic;
        D_reg_move_target: in     vl_logic;
        E_reg_move_target: in     vl_logic;
        Ci_reg_set      : in     vl_logic;
        NegA_reg_set    : in     vl_logic;
        A_reg_hi_set    : in     vl_logic;
        A_reg_lo_set    : in     vl_logic;
        B_reg_hi_set    : in     vl_logic;
        B_reg_lo_set    : in     vl_logic;
        C_reg_hi_set    : in     vl_logic;
        C_reg_lo_set    : in     vl_logic;
        A_reg_hi_clr    : in     vl_logic;
        A_reg_lo_clr    : in     vl_logic;
        B_reg_hi_clr    : in     vl_logic;
        B_reg_lo_clr    : in     vl_logic;
        C_reg_hi_clr    : in     vl_logic;
        C_reg_lo_clr    : in     vl_logic;
        move_from_ADC_RESULT_LSB: in     vl_logic;
        xfer_din_mux    : in     vl_logic_vector(31 downto 0);
        st_filt_curr_st : out    vl_logic;
        st_filt_next_qual: out    vl_logic;
        st_filt_0to1_eq : out    vl_logic;
        st_filt_1to0_eq : out    vl_logic;
        RRDIS2          : out    vl_logic;
        RRDIS1          : out    vl_logic;
        RRDIS0          : out    vl_logic;
        PPE_CTRL        : out    vl_logic_vector(31 downto 0);
        PPE_PC_ETC      : out    vl_logic_vector(31 downto 0);
        PPE_SCRATCH     : out    vl_logic_vector(31 downto 0);
        PPE_SF          : out    vl_logic_vector(31 downto 0);
        ALU_CTRL        : out    vl_logic_vector(31 downto 0);
        ALU_STATUS      : out    vl_logic_vector(31 downto 0);
        ALU_A           : out    vl_logic_vector(31 downto 0);
        ALU_B           : out    vl_logic_vector(31 downto 0);
        ALU_C           : out    vl_logic_vector(31 downto 0);
        ALU_D           : out    vl_logic_vector(15 downto 0);
        ALU_E           : out    vl_logic_vector(15 downto 0);
        C_reg_31        : out    vl_logic;
        PC_override     : out    vl_logic;
        PREADY_ALU      : out    vl_logic
    );
end F2DSS_ACE_PPE_ALU;
