library verilog;
use verilog.vl_types.all;
entity Matrix5x8 is
    port(
        HCLK            : in     vl_logic;
        HRESETn         : in     vl_logic;
        F2_TESTREMAPENABLE: in     vl_logic;
        F2_TESTESRAM1REMAP: in     vl_logic;
        F2_ESRAMSIZE    : in     vl_logic_vector(1 downto 0);
        F2_ENVMPOWEREDDOWN: in     vl_logic;
        COM_ESRAMFWREMAP: in     vl_logic;
        COM_ENVMREMAPSIZE: in     vl_logic_vector(4 downto 0);
        COM_ENVMREMAPBASE: in     vl_logic_vector(19 downto 0);
        COM_ENVMFABREMAPBASE: in     vl_logic_vector(19 downto 0);
        COM_PROTREGIONSIZE: in     vl_logic_vector(4 downto 0);
        COM_PROTREGIONBASE: in     vl_logic_vector(31 downto 0);
        COM_MASTERENABLE: in     vl_logic_vector(2 downto 0);
        COM_CLEARSTATUS : in     vl_logic_vector(4 downto 0);
        COM_WEIGHTEDMODE: in     vl_logic;
        COM_ERRORSTATUS : out    vl_logic_vector(4 downto 0);
        COM_ERRORINTERRUPT: out    vl_logic;
        HADDR_M0        : in     vl_logic_vector(31 downto 0);
        HMASTLOCK_M0    : in     vl_logic;
        HSIZE_M0        : in     vl_logic_vector(2 downto 0);
        HTRANS1_M0      : in     vl_logic;
        HWRITE_M0       : in     vl_logic;
        HWDATA_M0       : in     vl_logic_vector(31 downto 0);
        HRESP_M0        : out    vl_logic;
        HRDATA_M0       : out    vl_logic_vector(31 downto 0);
        HREADY_M0       : out    vl_logic;
        HADDR_M1        : in     vl_logic_vector(31 downto 0);
        HMASTLOCK_M1    : in     vl_logic;
        HSIZE_M1        : in     vl_logic_vector(2 downto 0);
        HTRANS1_M1      : in     vl_logic;
        HWRITE_M1       : in     vl_logic;
        HWDATA_M1       : in     vl_logic_vector(31 downto 0);
        HRESP_M1        : out    vl_logic;
        HRDATA_M1       : out    vl_logic_vector(31 downto 0);
        HREADY_M1       : out    vl_logic;
        HADDR_M2        : in     vl_logic_vector(31 downto 0);
        HMASTLOCK_M2    : in     vl_logic;
        HSIZE_M2        : in     vl_logic_vector(2 downto 0);
        HTRANS1_M2      : in     vl_logic;
        HWRITE_M2       : in     vl_logic;
        HWDATA_M2       : in     vl_logic_vector(31 downto 0);
        HRESP_M2        : out    vl_logic;
        HRDATA_M2       : out    vl_logic_vector(31 downto 0);
        HREADY_M2       : out    vl_logic;
        HADDR_M3        : in     vl_logic_vector(31 downto 0);
        HMASTLOCK_M3    : in     vl_logic;
        HSIZE_M3        : in     vl_logic_vector(2 downto 0);
        HTRANS1_M3      : in     vl_logic;
        HWRITE_M3       : in     vl_logic;
        HWDATA_M3       : in     vl_logic_vector(31 downto 0);
        HRESP_M3        : out    vl_logic;
        HRDATA_M3       : out    vl_logic_vector(31 downto 0);
        HREADY_M3       : out    vl_logic;
        HADDR_M4        : in     vl_logic_vector(31 downto 0);
        HMASTLOCK_M4    : in     vl_logic;
        HSIZE_M4        : in     vl_logic_vector(2 downto 0);
        HTRANS1_M4      : in     vl_logic;
        HWRITE_M4       : in     vl_logic;
        HWDATA_M4       : in     vl_logic_vector(31 downto 0);
        HRESP_M4        : out    vl_logic;
        HRDATA_M4       : out    vl_logic_vector(31 downto 0);
        HREADY_M4       : out    vl_logic;
        HRDATA_S0       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S0    : in     vl_logic;
        HRESP_S0        : in     vl_logic;
        HSEL_S0         : out    vl_logic;
        HADDR_S0        : out    vl_logic_vector(31 downto 0);
        HSIZE_S0        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S0      : out    vl_logic;
        HWRITE_S0       : out    vl_logic;
        HWDATA_S0       : out    vl_logic_vector(31 downto 0);
        HREADY_S0       : out    vl_logic;
        HRDATA_S1       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S1    : in     vl_logic;
        HRESP_S1        : in     vl_logic;
        HSEL_S1         : out    vl_logic;
        HADDR_S1        : out    vl_logic_vector(31 downto 0);
        HSIZE_S1        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S1      : out    vl_logic;
        HWRITE_S1       : out    vl_logic;
        HWDATA_S1       : out    vl_logic_vector(31 downto 0);
        HREADY_S1       : out    vl_logic;
        HRDATA_S2       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S2    : in     vl_logic;
        HRESP_S2        : in     vl_logic;
        HSEL_S2         : out    vl_logic;
        HADDR_S2        : out    vl_logic_vector(31 downto 0);
        HSIZE_S2        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S2      : out    vl_logic;
        HWRITE_S2       : out    vl_logic;
        HWDATA_S2       : out    vl_logic_vector(31 downto 0);
        HREADY_S2       : out    vl_logic;
        HRDATA_S3       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S3    : in     vl_logic;
        HRESP_S3        : in     vl_logic;
        HSEL_S3         : out    vl_logic;
        HADDR_S3        : out    vl_logic_vector(31 downto 0);
        HSIZE_S3        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S3      : out    vl_logic;
        HWRITE_S3       : out    vl_logic;
        HWDATA_S3       : out    vl_logic_vector(31 downto 0);
        HREADY_S3       : out    vl_logic;
        HRDATA_S4       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S4    : in     vl_logic;
        HRESP_S4        : in     vl_logic;
        HSEL_S4         : out    vl_logic;
        HADDR_S4        : out    vl_logic_vector(31 downto 0);
        HSIZE_S4        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S4      : out    vl_logic;
        HWRITE_S4       : out    vl_logic;
        HWDATA_S4       : out    vl_logic_vector(31 downto 0);
        HREADY_S4       : out    vl_logic;
        HRDATA_S5       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S5    : in     vl_logic;
        HRESP_S5        : in     vl_logic;
        HSEL_S5         : out    vl_logic;
        HADDR_S5        : out    vl_logic_vector(31 downto 0);
        HSIZE_S5        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S5      : out    vl_logic;
        HWRITE_S5       : out    vl_logic;
        HWDATA_S5       : out    vl_logic_vector(31 downto 0);
        HREADY_S5       : out    vl_logic;
        HMASTLOCK_S5    : out    vl_logic;
        HRDATA_S6       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S6    : in     vl_logic;
        HRESP_S6        : in     vl_logic;
        HSEL_S6         : out    vl_logic;
        HADDR_S6        : out    vl_logic_vector(31 downto 0);
        HSIZE_S6        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S6      : out    vl_logic;
        HWRITE_S6       : out    vl_logic;
        HWDATA_S6       : out    vl_logic_vector(31 downto 0);
        HREADY_S6       : out    vl_logic;
        HRDATA_S7       : in     vl_logic_vector(31 downto 0);
        HREADYOUT_S7    : in     vl_logic;
        HRESP_S7        : in     vl_logic;
        HSEL_S7         : out    vl_logic;
        HADDR_S7        : out    vl_logic_vector(31 downto 0);
        HSIZE_S7        : out    vl_logic_vector(2 downto 0);
        HTRANS1_S7      : out    vl_logic;
        HWRITE_S7       : out    vl_logic;
        HWDATA_S7       : out    vl_logic_vector(31 downto 0);
        HREADY_S7       : out    vl_logic
    );
end Matrix5x8;
