----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Oct 19 12:51:53 2011
-- Testbench Template
-- This is a basic testbench that instantiates your design with basic 
-- clock and reset pins connected.  If your design has special
-- clock/reset or testbench driver requirements then you should 
-- copy this file and modify it. 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity testbench is
end testbench;

architecture behavioral of testbench is

    constant SYSCLK_PERIOD : time := 100 ns;

    signal SYSCLK : std_logic := '0';
    signal NSYSRESET : std_logic := '0';

    component complex_mult
        -- ports
        port( 
            -- Inputs
            sample_rdy_in : in std_logic;
            CLK : in std_logic;
            RST : in std_logic;
            I_A : in std_logic_vector(7 downto 0);
            I_B : in std_logic_vector(13 downto 0);
            Q_A : in std_logic_vector(7 downto 0);
            Q_B : in std_logic_vector(13 downto 0);

            -- Outputs
            I : out std_logic_vector(22 downto 0);
            Q : out std_logic_vector(22 downto 0)

            -- Inouts

        );
    end component;

begin

    process
        variable vhdl_initial : BOOLEAN := TRUE;

    begin
        if ( vhdl_initial ) then
            -- Assert Reset
            NSYSRESET <= '0';
            wait for ( SYSCLK_PERIOD * 10 );
            
            NSYSRESET <= '1';
            wait;
        end if;
    end process;

    -- 10MHz Clock Driver
    SYSCLK <= not SYSCLK after (SYSCLK_PERIOD / 2.0 );

    -- Instantiate Unit Under Test:  complex_mult
    complex_mult_0 : complex_mult
        -- port map
        port map( 
            -- Inputs
            sample_rdy_in => '0',
            CLK => SYSCLK,
            RST => NSYSRESET,
            I_A => (others=> '0'),
            I_B => (others=> '0'),
            Q_A => (others=> '0'),
            Q_B => (others=> '0'),

            -- Outputs
            I => open,
            Q => open

            -- Inouts

        );

end behavioral;

