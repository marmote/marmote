----------------------------------------------------------------------
-- Created by Actel SmartDesign Wed Nov 23 15:32:40 2011
-- Testbench Template
-- This is a basic testbench that instantiates your design with basic 
-- clock and reset pins connected.  If your design has special
-- clock/reset or testbench driver requirements then you should 
-- copy this file and modify it. 
----------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity testbench is
end testbench;

architecture behavioral of testbench is

    constant SYSCLK_PERIOD : time := 100 ns;

    signal SYSCLK : std_logic := '0';
    signal NSYSRESET : std_logic := '0';

    component DDC
        -- ports
        port( 
            -- Inputs
            RST : in std_logic;
            CLK : in std_logic;
            sample_rdy_in : in std_logic;
            I_in : in std_logic_vector(13 downto 0);
            Q_in : in std_logic_vector(13 downto 0);
            DPHASE : in std_logic_vector(15 downto 0);
            I_DC_cor : in std_logic_vector(13 downto 0);
            Q_DC_cor : in std_logic_vector(13 downto 0);

            -- Outputs
            I_SMPL_RDY : out std_logic;
            Q_SMPL_RDY : out std_logic;
            I_out : out std_logic_vector(26 downto 0);
            Q_out : out std_logic_vector(26 downto 0)

            -- Inouts

        );
    end component;

begin

    process
        variable vhdl_initial : BOOLEAN := TRUE;

    begin
        if ( vhdl_initial ) then
            -- Assert Reset
            NSYSRESET <= '0';
            wait for ( SYSCLK_PERIOD * 10 );
            
            NSYSRESET <= '1';
            wait;
        end if;
    end process;

    -- 10MHz Clock Driver
    SYSCLK <= not SYSCLK after (SYSCLK_PERIOD / 2.0 );

    -- Instantiate Unit Under Test:  DDC
    DDC_0 : DDC
        -- port map
        port map( 
            -- Inputs
            RST => NSYSRESET,
            CLK => SYSCLK,
            sample_rdy_in => '0',
            I_in => (others=> '0'),
            Q_in => (others=> '0'),
            DPHASE => (others=> '0'),
            I_DC_cor => (others=> '0'),
            Q_DC_cor => (others=> '0'),

            -- Outputs
            I_SMPL_RDY =>  open,
            Q_SMPL_RDY =>  open,
            I_out => open,
            Q_out => open

            -- Inouts

        );

end behavioral;

