----------------------------------------------------------------------
-- Created by Actel SmartDesign Tue Jul 19 15:02:10 2011
-- Parameters for CORECORDIC
----------------------------------------------------------------------


package coreparameters is
    constant ARCH : integer := 1;
    constant BIT_WIDTH : integer := 16;
    constant FAMILY : integer := 15;
    constant HDL_license : string( 1 to 1 ) := "U";
    constant ITERATIONS : integer := 16;
    constant MODE : integer := 0;
    constant testbench : string( 1 to 4 ) := "User";
end coreparameters;
