library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_PPE is
    port(
        PCLK            : in     vl_logic;
        PRESETN         : in     vl_logic;
        PADDR           : in     vl_logic_vector(12 downto 0);
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PRDATA_PPE      : out    vl_logic_vector(31 downto 0);
        PREADY_PPE      : out    vl_logic;
        PPE2SSE_PSEL    : out    vl_logic;
        PPE2SSE_PENABLE : out    vl_logic;
        PPE2SSE_PWRITE  : out    vl_logic;
        PPE2SSE_PADDR   : out    vl_logic_vector(11 downto 0);
        PPE2SSE_PWDATA  : out    vl_logic_vector(15 downto 0);
        PPE2SSE_PRDATA  : in     vl_logic_vector(15 downto 0);
        PPE2SSE_PREADY  : in     vl_logic;
        PPE2SSE_STALL   : out    vl_logic;
        PPE_BUSY        : out    vl_logic;
        SSE_ADC0_RESULTS: in     vl_logic;
        SSE_ADC1_RESULTS: in     vl_logic;
        SSE_ADC2_RESULTS: in     vl_logic;
        ADC0_DATAVALID_rise: in     vl_logic;
        ADC1_DATAVALID_rise: in     vl_logic;
        ADC2_DATAVALID_rise: in     vl_logic;
        ADC0_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC1_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC2_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC0_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC1_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC2_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        PPE_FLAGS0      : out    vl_logic_vector(31 downto 0);
        PPE_FLAGS1      : out    vl_logic_vector(31 downto 0);
        PPE_FLAGS2      : out    vl_logic_vector(31 downto 0);
        PPE_FLAGS3      : out    vl_logic_vector(31 downto 0);
        PPE_SFFLAGS     : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_FULL  : out    vl_logic;
        ADC0_FIFO_AFULL : out    vl_logic;
        ADC1_FIFO_FULL  : out    vl_logic;
        ADC1_FIFO_AFULL : out    vl_logic;
        ADC2_FIFO_FULL  : out    vl_logic;
        ADC2_FIFO_AFULL : out    vl_logic;
        ADC0_FIFO_EMPTY : out    vl_logic;
        ADC1_FIFO_EMPTY : out    vl_logic;
        ADC2_FIFO_EMPTY : out    vl_logic;
        PPE_PDMA_DATAOUT_reg_move_target: out    vl_logic;
        PPE_PDMA_DATAOUT_chan_en: out    vl_logic;
        PPE_PDMA_DATAOUT_raw_en: out    vl_logic;
        PPE_PDMA_DATAOUT_tag_en: out    vl_logic;
        PPE_PDMA_CTRL_reg_move_target: out    vl_logic;
        xfer_din_mux    : out    vl_logic_vector(31 downto 0);
        CURRENT_ADC_CHAN: out    vl_logic_vector(5 downto 0);
        TEST_MODE       : in     vl_logic;
        RB_TEST         : in     vl_logic;
        RB_CSBA         : in     vl_logic;
        RB_CSBB         : in     vl_logic;
        RB_RWBA         : in     vl_logic;
        RB_RWBB         : in     vl_logic;
        RB_ADA          : in     vl_logic_vector(8 downto 0);
        RB_ADB          : in     vl_logic_vector(8 downto 0);
        RB_WDA          : in     vl_logic_vector(31 downto 0);
        RB_WDB          : in     vl_logic_vector(31 downto 0);
        RB_RDA          : out    vl_logic_vector(31 downto 0);
        RB_RDB          : out    vl_logic_vector(31 downto 0)
    );
end F2DSS_ACE_PPE;
