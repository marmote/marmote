----------------------------------------------------------------------
-- Created by Actel SmartDesign Thu May 26 11:49:35 2011
-- Parameters for CORESPI
----------------------------------------------------------------------


package coreparameters is
    constant FAMILY : integer := 15;
    constant HDL_license : string( 1 to 1 ) := "O";
    constant testbench : string( 1 to 4 ) := "User";
    constant USE_MASTER : integer := 1;
    constant USE_SLAVE : integer := 0;
end coreparameters;
