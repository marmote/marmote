library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_PPE_FIFO_CTRL is
    port(
        PCLK            : in     vl_logic;
        PRESETN         : in     vl_logic;
        PADDR           : in     vl_logic_vector(12 downto 0);
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PREADY_FIFO_CTRL: out    vl_logic;
        xfer_din_mux    : in     vl_logic_vector(31 downto 0);
        PPE2SSE_PSEL    : in     vl_logic;
        PPE2SSE_PWDATA  : in     vl_logic_vector(15 downto 0);
        PPE2SSE_STALL   : out    vl_logic;
        ADC_FIFO_rd     : in     vl_logic;
        ADC0_FIFO_CTRL_reg_move_target: in     vl_logic;
        ADC1_FIFO_CTRL_reg_move_target: in     vl_logic;
        ADC2_FIFO_CTRL_reg_move_target: in     vl_logic;
        SSE_ADC0_RESULTS: in     vl_logic;
        SSE_ADC1_RESULTS: in     vl_logic;
        SSE_ADC2_RESULTS: in     vl_logic;
        ADC0_DATAVALID_rise: in     vl_logic;
        ADC1_DATAVALID_rise: in     vl_logic;
        ADC2_DATAVALID_rise: in     vl_logic;
        ADC0_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC1_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC2_RESULT     : in     vl_logic_vector(11 downto 0);
        ADC0_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC1_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC2_CHNUMBER   : in     vl_logic_vector(4 downto 0);
        ADC_FIFO_PTR_inc: in     vl_logic;
        ADC_FIFO_PTR_clr: in     vl_logic;
        ADC_FIFO_PTR    : out    vl_logic_vector(1 downto 0);
        RAM_DO_B        : in     vl_logic_vector(31 downto 0);
        PC_init_addr    : out    vl_logic_vector(9 downto 0);
        CURRENT_ADC_CHAN: out    vl_logic_vector(5 downto 0);
        CURRENT_ADC_RESULT: out    vl_logic_vector(11 downto 0);
        ADC0_FIFO_FULL  : out    vl_logic;
        ADC0_FIFO_AFULL : out    vl_logic;
        ADC1_FIFO_FULL  : out    vl_logic;
        ADC1_FIFO_AFULL : out    vl_logic;
        ADC2_FIFO_FULL  : out    vl_logic;
        ADC2_FIFO_AFULL : out    vl_logic;
        ADC0_FIFO_EMPTY : out    vl_logic;
        ADC1_FIFO_EMPTY : out    vl_logic;
        ADC2_FIFO_EMPTY : out    vl_logic;
        ADC_FIFO_EMPTY  : out    vl_logic;
        OTHER_ADC_FIFOS_NOT_EMPTY: out    vl_logic;
        RRDIS0          : in     vl_logic;
        RRDIS1          : in     vl_logic;
        RRDIS2          : in     vl_logic;
        RR_DISABLE      : out    vl_logic;
        ADC0_FIFO_CTRL  : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_STATUS: out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA  : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA_PEEK: out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA0 : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA1 : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA2 : out    vl_logic_vector(31 downto 0);
        ADC0_FIFO_DATA3 : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_CTRL  : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_STATUS: out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA  : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA_PEEK: out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA0 : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA1 : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA2 : out    vl_logic_vector(31 downto 0);
        ADC1_FIFO_DATA3 : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_CTRL  : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_STATUS: out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA  : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA_PEEK: out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA0 : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA1 : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA2 : out    vl_logic_vector(31 downto 0);
        ADC2_FIFO_DATA3 : out    vl_logic_vector(31 downto 0)
    );
end F2DSS_ACE_PPE_FIFO_CTRL;
