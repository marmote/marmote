library verilog;
use verilog.vl_types.all;
entity F2DSS_ACE_PPE_FSM is
    port(
        PCLK            : in     vl_logic;
        PRESETN         : in     vl_logic;
        PC_override     : in     vl_logic;
        PPE_CTRL        : in     vl_logic_vector(31 downto 0);
        PPE_PC_ETC      : in     vl_logic_vector(31 downto 0);
        PPE_FPTR        : in     vl_logic_vector(31 downto 0);
        RAM_DO_A        : in     vl_logic_vector(31 downto 0);
        RAM_ADDRESSES_EQUAL: in     vl_logic;
        RAM_RD_A        : out    vl_logic;
        RAM_RD_B        : out    vl_logic;
        RAM_RD_B_hold_en: out    vl_logic;
        RAM_WR_B        : out    vl_logic;
        RAM_ADDR_A      : out    vl_logic_vector(8 downto 0);
        RAM_ADDR_B      : out    vl_logic_vector(8 downto 0);
        PPE_BUSY        : out    vl_logic;
        PPE2SSE_PREADY  : in     vl_logic;
        PPE2SSE_wr      : out    vl_logic;
        PPE2SSE_rd_hold_en: out    vl_logic;
        PPE2SSE_sel     : out    vl_logic;
        PPE2SSE_en      : out    vl_logic;
        st_filt_curr_st : in     vl_logic;
        st_filt_next_qual: in     vl_logic;
        st_filt_0to1_eq : in     vl_logic;
        st_filt_1to0_eq : in     vl_logic;
        C_reg_31        : in     vl_logic;
        CURRENT_ADC_CHAN: in     vl_logic_vector(5 downto 0);
        ADC_FIFO_EMPTY  : in     vl_logic;
        OTHER_ADC_FIFOS_NOT_EMPTY: in     vl_logic;
        RR_DISABLE      : in     vl_logic;
        ADC_FIFO_PTR_inc: out    vl_logic;
        ADC_FIFO_PTR_clr: out    vl_logic;
        ADC_FIFO_rd     : out    vl_logic;
        ADC0_FIFO_CTRL_reg_move_target: out    vl_logic;
        ADC1_FIFO_CTRL_reg_move_target: out    vl_logic;
        ADC2_FIFO_CTRL_reg_move_target: out    vl_logic;
        st_filt_cnt_clr : out    vl_logic;
        st_filt_cnt_inc : out    vl_logic;
        st_filt_st_one  : out    vl_logic;
        st_filt_st_zero : out    vl_logic;
        PC_init_addr_ld : out    vl_logic;
        PC_inc          : out    vl_logic;
        PC_ETC_busy     : out    vl_logic;
        SF_busy         : out    vl_logic;
        THR_busy        : out    vl_logic;
        SCRATCH_busy    : out    vl_logic;
        ALU_CTRL_busy   : out    vl_logic;
        A_busy          : out    vl_logic;
        B_busy          : out    vl_logic;
        C_busy          : out    vl_logic;
        D_busy          : out    vl_logic;
        E_busy          : out    vl_logic;
        Ci_busy         : out    vl_logic;
        NegA_busy       : out    vl_logic;
        C2a_busy        : out    vl_logic;
        s2B_busy        : out    vl_logic;
        C2d_busy        : out    vl_logic;
        PPE_FPTR_busy   : out    vl_logic;
        PPE_FLAGS0_busy : out    vl_logic;
        PPE_FLAGS1_busy : out    vl_logic;
        PPE_FLAGS2_busy : out    vl_logic;
        PPE_FLAGS3_busy : out    vl_logic;
        PPE_SFFLAGS_busy: out    vl_logic;
        xfer_load_special_active: out    vl_logic;
        xfer_move_active: out    vl_logic;
        PPE_CTRL_reg_move_target: out    vl_logic;
        PC_ETC_reg_move_target: out    vl_logic;
        SCRATCH_reg_move_target: out    vl_logic;
        SF_reg_move_target: out    vl_logic;
        ALU_CTRL_reg_move_target: out    vl_logic;
        A_reg_move_target: out    vl_logic;
        B_reg_move_target: out    vl_logic;
        C_reg_move_target: out    vl_logic;
        D_reg_move_target: out    vl_logic;
        E_reg_move_target: out    vl_logic;
        PPE_FPTR_reg_move_target: out    vl_logic;
        PPE_FLAGS0_reg_move_target: out    vl_logic;
        PPE_FLAGS1_reg_move_target: out    vl_logic;
        PPE_FLAGS2_reg_move_target: out    vl_logic;
        PPE_FLAGS3_reg_move_target: out    vl_logic;
        PPE_SFFLAGS_reg_move_target: out    vl_logic;
        PPE2SSE_PADDR_reg_move_target: out    vl_logic;
        PPE2SSE_PWDATA_LSB_reg_move_target: out    vl_logic;
        PPE2SSE_PWDATA_MSB_reg_move_target: out    vl_logic;
        PPE_PDMA_DATAOUT_reg_move_target: out    vl_logic;
        PPE_PDMA_DATAOUT_chan_en: out    vl_logic;
        PPE_PDMA_DATAOUT_raw_en: out    vl_logic;
        PPE_PDMA_DATAOUT_tag_en: out    vl_logic;
        PPE_PDMA_CTRL_reg_move_target: out    vl_logic;
        PPE_FLAG_bit    : out    vl_logic;
        PPE_FLAG_bit_update: out    vl_logic;
        PPE_thresh_op_load: out    vl_logic;
        move_from_PPE_CTRL: out    vl_logic;
        move_from_PC_ETC: out    vl_logic;
        move_from_SF    : out    vl_logic;
        move_from_SCRATCH: out    vl_logic;
        move_from_ALU_CTRL: out    vl_logic;
        move_from_ALU_STATUS: out    vl_logic;
        move_from_A     : out    vl_logic;
        move_from_B     : out    vl_logic;
        move_from_C     : out    vl_logic;
        move_from_PPE_FPTR: out    vl_logic;
        move_from_PPE_FLAGS0: out    vl_logic;
        move_from_PPE_FLAGS1: out    vl_logic;
        move_from_PPE_FLAGS2: out    vl_logic;
        move_from_PPE_FLAGS3: out    vl_logic;
        move_from_PPE_SFFLAGS: out    vl_logic;
        move_from_ADC0_FIFO_CTRL: out    vl_logic;
        move_from_ADC0_FIFO_STATUS: out    vl_logic;
        move_from_ADC0_FIFO_DATA: out    vl_logic;
        move_from_ADC1_FIFO_CTRL: out    vl_logic;
        move_from_ADC1_FIFO_STATUS: out    vl_logic;
        move_from_ADC1_FIFO_DATA: out    vl_logic;
        move_from_ADC2_FIFO_CTRL: out    vl_logic;
        move_from_ADC2_FIFO_STATUS: out    vl_logic;
        move_from_ADC2_FIFO_DATA: out    vl_logic;
        move_from_ADC_RESULT_LSB: out    vl_logic;
        move_from_ADC_RESULT_MSB: out    vl_logic;
        move_from_PPE2SSE_PRDATA: out    vl_logic;
        move_from_RAM_DO_A_31_0: out    vl_logic;
        move_from_RAM_DO_A_23_0_LSB: out    vl_logic;
        move_from_RAM_DO_A_23_0_MSB: out    vl_logic;
        move_from_RAM_DO_A_15_0_MSB: out    vl_logic;
        move_from_RAM_DO_B_31_0: out    vl_logic;
        RAM_DI_B_31_0_move_target: out    vl_logic;
        RAM_DI_B_23_0_move_target: out    vl_logic;
        RAM_DI_B_15_0_move_target: out    vl_logic;
        keep_bits_31_24 : out    vl_logic;
        keep_bits_7_0   : out    vl_logic;
        Ci_reg_set      : out    vl_logic;
        NegA_reg_set    : out    vl_logic;
        A_reg_hi_set    : out    vl_logic;
        A_reg_lo_set    : out    vl_logic;
        B_reg_hi_set    : out    vl_logic;
        B_reg_lo_set    : out    vl_logic;
        C_reg_hi_set    : out    vl_logic;
        C_reg_lo_set    : out    vl_logic;
        A_reg_hi_clr    : out    vl_logic;
        A_reg_lo_clr    : out    vl_logic;
        B_reg_hi_clr    : out    vl_logic;
        B_reg_lo_clr    : out    vl_logic;
        C_reg_hi_clr    : out    vl_logic;
        C_reg_lo_clr    : out    vl_logic
    );
end F2DSS_ACE_PPE_FSM;
