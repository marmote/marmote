library verilog;
use verilog.vl_types.all;
entity F2DSS_SSE is
    port(
        PRESETN         : in     vl_logic;
        PCLK            : in     vl_logic;
        HCLK            : in     vl_logic;
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PWRITE          : in     vl_logic;
        PADDR           : in     vl_logic_vector(11 downto 0);
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PRDATA          : out    vl_logic_vector(15 downto 0);
        PREADY          : out    vl_logic;
        PSLVERR         : out    vl_logic;
        PPE_PSEL        : in     vl_logic;
        PPE_PENABLE     : in     vl_logic;
        PPE_PWRITE      : in     vl_logic;
        PPE_PADDR       : in     vl_logic_vector(11 downto 0);
        PPE_PWDATA      : in     vl_logic_vector(15 downto 0);
        PPE_PRDATA      : out    vl_logic_vector(15 downto 0);
        PPE_PREADY      : out    vl_logic;
        PPE_PSLVERR     : out    vl_logic;
        PPE_FIFO_FULL   : in     vl_logic;
        PC0_FLAGS       : out    vl_logic_vector(3 downto 0);
        PC1_FLAGS       : out    vl_logic_vector(3 downto 0);
        PC2_FLAGS       : out    vl_logic_vector(3 downto 0);
        ADC0_CALIBRATE_rise: out    vl_logic;
        ADC1_CALIBRATE_rise: out    vl_logic;
        ADC2_CALIBRATE_rise: out    vl_logic;
        ADC0_CALIBRATE_fall: out    vl_logic;
        ADC1_CALIBRATE_fall: out    vl_logic;
        ADC2_CALIBRATE_fall: out    vl_logic;
        ADC0_DATAVALID_rise: out    vl_logic;
        ADC1_DATAVALID_rise: out    vl_logic;
        ADC2_DATAVALID_rise: out    vl_logic;
        FPGA_TRIGGER    : in     vl_logic;
        ADC0_BUSY       : in     vl_logic;
        ADC1_BUSY       : in     vl_logic;
        ADC2_BUSY       : in     vl_logic;
        ADC0_CALIBRATE  : in     vl_logic;
        ADC1_CALIBRATE  : in     vl_logic;
        ADC2_CALIBRATE  : in     vl_logic;
        ADC0_DATAVALID  : in     vl_logic;
        ADC1_DATAVALID  : in     vl_logic;
        ADC2_DATAVALID  : in     vl_logic;
        ADC0_SAMPLE     : in     vl_logic;
        ADC1_SAMPLE     : in     vl_logic;
        ADC2_SAMPLE     : in     vl_logic;
        ADC0_TVC        : out    vl_logic_vector(7 downto 0);
        ADC1_TVC        : out    vl_logic_vector(7 downto 0);
        ADC2_TVC        : out    vl_logic_vector(7 downto 0);
        ADC0_STC        : out    vl_logic_vector(7 downto 0);
        ADC1_STC        : out    vl_logic_vector(7 downto 0);
        ADC2_STC        : out    vl_logic_vector(7 downto 0);
        ADC0_MODE       : out    vl_logic_vector(3 downto 0);
        ADC1_MODE       : out    vl_logic_vector(3 downto 0);
        ADC2_MODE       : out    vl_logic_vector(3 downto 0);
        ADC_VAREFSEL    : out    vl_logic;
        ABPOWERON       : out    vl_logic;
        ADC0_CHNUMBER   : out    vl_logic_vector(4 downto 0);
        ADC1_CHNUMBER   : out    vl_logic_vector(4 downto 0);
        ADC2_CHNUMBER   : out    vl_logic_vector(4 downto 0);
        ADC0_ADCSTART   : out    vl_logic;
        ADC1_ADCSTART   : out    vl_logic;
        ADC2_ADCSTART   : out    vl_logic;
        ADC0_PWRDWN     : out    vl_logic;
        ADC1_PWRDWN     : out    vl_logic;
        ADC2_PWRDWN     : out    vl_logic;
        ADC0_ADCRESET   : out    vl_logic;
        ADC1_ADCRESET   : out    vl_logic;
        ADC2_ADCRESET   : out    vl_logic;
        ACB_RDATA       : in     vl_logic_vector(7 downto 0);
        ACB_ADDR        : out    vl_logic_vector(7 downto 0);
        ACB_WRE         : out    vl_logic;
        ACB_WDATA       : out    vl_logic_vector(7 downto 0);
        ACB_RESETN      : out    vl_logic;
        OBD_FPGA0_CLKOUT: in     vl_logic;
        OBD_FPGA1_CLKOUT: in     vl_logic;
        OBD_FPGA2_CLKOUT: in     vl_logic;
        OBD_FPGA0_DOUT  : in     vl_logic;
        OBD_FPGA1_DOUT  : in     vl_logic;
        OBD_FPGA2_DOUT  : in     vl_logic;
        OBD_DOUT0       : out    vl_logic;
        OBD_DOUT1       : out    vl_logic;
        OBD_DOUT2       : out    vl_logic;
        OBD_CLKOUT0     : out    vl_logic;
        OBD_CLKOUT1     : out    vl_logic;
        OBD_CLKOUT2     : out    vl_logic;
        OBD_ENABLE0     : out    vl_logic;
        OBD_ENABLE1     : out    vl_logic;
        OBD_ENABLE2     : out    vl_logic;
        INREADY         : out    vl_logic;
        SSE_ADC0_RESULTS: out    vl_logic;
        SSE_ADC1_RESULTS: out    vl_logic;
        SSE_ADC2_RESULTS: out    vl_logic
    );
end F2DSS_SSE;
